 ----------------------------------------------------------------------------------
-- Company: Tu Delft
-- Engineer: HS Jagadeeshwar
-- 
-- Create Date: 10/02/2017 05:06:32 PM
-- Design Name: StimG_v1_4
-- Module Name: StimG_v1_4 - Behavioral
-- Project Name: Stimulus Generator
-- Target Devices: Zybo 
-- Tool Versions: Vivado 2015.4
-- Description: Top level module with component instantiation 
-- Dependencies: StimG_v1_4_S00_AXI and top 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments: Uses autogenerated templet from Xilinx IP packager after editing 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity StimG_v1_4 is
	generic (
		-- Users to add parameters here
        pulse_number : INTEGER := 4;
        pulse_number_bits : INTEGER := 2;
        PhyC : INTEGER := 2;
        StimC : INTEGER := 10;
        StimC_bits : INTEGER := 4;
        Clock_div : INTEGER := 5000;
        FIFO_size : INTEGER := 1024;
		-- User parameters ends
		-- Do not modify the parameters beyond this line
		-- Parameters of Axi Slave Bus Interface S00_AXI
		C_S00_AXI_DATA_WIDTH	: integer	:= 32;
		C_S00_AXI_ADDR_WIDTH	: integer	:= 5
	);
	port (
		-- Users to add ports here         
        M_AXIS_ACLK    : in std_logic;
        M_AXIS_ARESETN : in std_logic;
        cluster_rdy    : in STD_LOGIC;
        cluster_in_ack : in STD_LOGIC;
        cluster_in_str : out STD_LOGIC;
        cluster_in_type : out STD_LOGIC_VECTOR (1 downto 0);
        cluster_in_data : out STD_LOGIC_VECTOR (31 downto 0);
        cluster_in_adr : out STD_LOGIC_VECTOR (StimC_bits-1 downto 0);   
		-- User ports ends
		-- Do not modify the ports beyond this line


		-- Ports of Axi Slave Bus Interface S00_AXI
		s00_axi_aclk	: in std_logic;
		s00_axi_aresetn	: in std_logic;
		s00_axi_awaddr	: in std_logic_vector(C_S00_AXI_ADDR_WIDTH-1 downto 0);
		s00_axi_awprot	: in std_logic_vector(2 downto 0);
		s00_axi_awvalid	: in std_logic;
		s00_axi_awready	: out std_logic;
		s00_axi_wdata	: in std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
		s00_axi_wstrb	: in std_logic_vector((C_S00_AXI_DATA_WIDTH/8)-1 downto 0);
		s00_axi_wvalid	: in std_logic;
		s00_axi_wready	: out std_logic;
		s00_axi_bresp	: out std_logic_vector(1 downto 0);
		s00_axi_bvalid	: out std_logic;
		s00_axi_bready	: in std_logic;
		s00_axi_araddr	: in std_logic_vector(C_S00_AXI_ADDR_WIDTH-1 downto 0);
		s00_axi_arprot	: in std_logic_vector(2 downto 0);
		s00_axi_arvalid	: in std_logic;
		s00_axi_arready	: out std_logic;
		s00_axi_rdata	: out std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
		s00_axi_rresp	: out std_logic_vector(1 downto 0);
		s00_axi_rvalid	: out std_logic;
		s00_axi_rready	: in std_logic
	);
end StimG_v1_4;

architecture arch_imp of StimG_v1_4 is

	-- component declaration
	component StimG_v1_4_S00_AXI is
		generic (
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		C_S_AXI_ADDR_WIDTH	: integer	:= 5;
			 StimC_bits : INTEGER := 4;
            pulse_number_bits : INTEGER := 2
		);
		port (
				start         : OUT STD_LOGIC;
        init_str    : OUT STD_LOGIC;
        init_in_typ    : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        cell_in_address : OUT STD_LOGIC_VECTOR(StimC_bits-1 DOWNTO 0) ;
        pulse_in_address: OUT  STD_LOGIC_VECTOR(pulse_number_bits-1 DOWNTO 0);
        init_in_data_top: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        init_ack    : IN STD_LOGIC;
        start_ack    : IN STD_LOGIC;
		S_AXI_ACLK	: in std_logic;
		S_AXI_ARESETN	: in std_logic;
		S_AXI_AWADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		S_AXI_AWPROT	: in std_logic_vector(2 downto 0);
		S_AXI_AWVALID	: in std_logic;
		S_AXI_AWREADY	: out std_logic;
		S_AXI_WDATA	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_WSTRB	: in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		S_AXI_WVALID	: in std_logic;
		S_AXI_WREADY	: out std_logic;
		S_AXI_BRESP	: out std_logic_vector(1 downto 0);
		S_AXI_BVALID	: out std_logic;
		S_AXI_BREADY	: in std_logic;
		S_AXI_ARADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		S_AXI_ARPROT	: in std_logic_vector(2 downto 0);
		S_AXI_ARVALID	: in std_logic;
		S_AXI_ARREADY	: out std_logic;
		S_AXI_RDATA	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_RRESP	: out std_logic_vector(1 downto 0);
		S_AXI_RVALID	: out std_logic;
		S_AXI_RREADY	: in std_logic
		);
	end component StimG_v1_4_S00_AXI;
		-----------------------------------------------------------------------------------------------------------------
        COMPONENT top IS
        -----------------------------------------------------------------------------------------------------------------
	    GENERIC (
        pulse_number : INTEGER := 4;
        pulse_number_bits : INTEGER := 2;
        PhyC : INTEGER := 2;
        StimC : INTEGER := 10;
        StimC_bits : INTEGER := 4;
        Clock_div : INTEGER := 2500;
        FIFO_size : INTEGER := 1024
    );
     port (
                M_AXIS_ACLK    : in std_logic;
                M_AXIS_ARESETN : in std_logic;
                cluster_rdy    : in STD_LOGIC;
                cluster_in_ack : in STD_LOGIC;
                cluster_in_str : out STD_LOGIC;
                cluster_in_type : out STD_LOGIC_VECTOR (1 downto 0);
                cluster_in_data : out STD_LOGIC_VECTOR (31 downto 0);
                cluster_in_adr : out STD_LOGIC_VECTOR (StimC_bits-1 downto 0);
                reset         : IN STD_LOGIC;
                clock         : IN STD_LOGIC;
                start         : IN STD_LOGIC;
                init_str    : IN STD_LOGIC;
                init_in_typ    : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
                cell_in_address : IN STD_LOGIC_VECTOR(StimC_bits-1 DOWNTO 0) ;
                pulse_in_address: IN  STD_LOGIC_VECTOR(pulse_number_bits-1 DOWNTO 0);
                init_in_data_top: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
                init_ack    : OUT STD_LOGIC;   
                start_ack    : OUT STD_LOGIC
     );
    END COMPONENT top;
	SIGNAL start         : STD_LOGIC;
    SIGNAL init_str    : STD_LOGIC;
    SIGNAL init_in_typ    :  STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL cell_in_address :  STD_LOGIC_VECTOR(StimC_bits-1 DOWNTO 0) ;
    SIGNAL pulse_in_address:   STD_LOGIC_VECTOR(pulse_number_bits-1 DOWNTO 0);
    SIGNAL init_in_data_top:  STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL init_ack    :  STD_LOGIC;
    SIGNAL start_ack   :  STD_LOGIC;
begin

-- Instantiation of Axi Bus Interface S00_AXI
StimG_v1_4_S00_AXI_inst : StimG_v1_4_S00_AXI
	generic map (
		C_S_AXI_DATA_WIDTH	=> C_S00_AXI_DATA_WIDTH,
		C_S_AXI_ADDR_WIDTH	=> C_S00_AXI_ADDR_WIDTH,
		StimC_bits => StimC_bits,
                pulse_number_bits => pulse_number_bits)
	port map (
		start=> start,
        init_str => init_str,
        init_in_typ => init_in_typ,  
        cell_in_address => cell_in_address,
        pulse_in_address => pulse_in_address,
        init_in_data_top => init_in_data_top,
        init_ack   => init_ack,
        start_ack  => start_ack,
		S_AXI_ACLK	=> s00_axi_aclk,
		S_AXI_ARESETN	=> s00_axi_aresetn,
		S_AXI_AWADDR	=> s00_axi_awaddr,
		S_AXI_AWPROT	=> s00_axi_awprot,
		S_AXI_AWVALID	=> s00_axi_awvalid,
		S_AXI_AWREADY	=> s00_axi_awready,
		S_AXI_WDATA	=> s00_axi_wdata,
		S_AXI_WSTRB	=> s00_axi_wstrb,
		S_AXI_WVALID	=> s00_axi_wvalid,
		S_AXI_WREADY	=> s00_axi_wready,
		S_AXI_BRESP	=> s00_axi_bresp,
		S_AXI_BVALID	=> s00_axi_bvalid,
		S_AXI_BREADY	=> s00_axi_bready,
		S_AXI_ARADDR	=> s00_axi_araddr,
		S_AXI_ARPROT	=> s00_axi_arprot,
		S_AXI_ARVALID	=> s00_axi_arvalid,
		S_AXI_ARREADY	=> s00_axi_arready,
		S_AXI_RDATA	=> s00_axi_rdata,
		S_AXI_RRESP	=> s00_axi_rresp,
		S_AXI_RVALID	=> s00_axi_rvalid,
		S_AXI_RREADY	=> s00_axi_rready
	);

	-- Add user logic here
uut_top : COMPONENT top
            GENERIC MAP (
            pulse_number,
            pulse_number_bits ,
            PhyC ,
            StimC ,
            StimC_bits,
            Clock_div,
            FIFO_size
           )
            PORT MAP(     
                    M_AXIS_ACLK => M_AXIS_ACLK,
                    M_AXIS_ARESETN => M_AXIS_ARESETN,
                    cluster_rdy => cluster_rdy,
                    cluster_in_ack => cluster_in_ack,
                    cluster_in_str => cluster_in_str,
                    cluster_in_type => cluster_in_type,
                    cluster_in_data => cluster_in_data,
                    cluster_in_adr => cluster_in_adr,
                    reset => M_AXIS_ARESETN, 
                    clock => M_AXIS_ACLK,
                    start=> start,
                    init_str => init_str, 
                    init_in_typ => init_in_typ, 
                    cell_in_address => cell_in_address, 
                    pulse_in_address => pulse_in_address, 
                    init_in_data_top => init_in_data_top, 
                    init_ack => init_ack,
                    start_ack => start_ack
            );
	-- User logic ends

end arch_imp;
